// wallace tb
module wallace_tb;

logic [31:0] a;
logic [31:0] b;
logic [63:0] s;
wallace w (
  .a(a), .b(b), .s(s)
);

initial begin
  #200ns;
  a <= 32'b11111111111111111111111111111111;
  b <= 32'b11111111111111111111111111111111;
  #20000ns;
  a <= 32'b00000000000000000000000000000000;
  b <= 32'b00000000000000000000000000000000;
  #20000ns;
  a <= 32'b00000000000000001001000100101001;
  b <= 32'b00000000000000001001000100010001;
  #20000ns;
end

endmodule

/*
a = 00000000000000001001000100101001
b = 00000000000000001001000100010001

row 1 should be 
  00000000000000001001000100101001
 00000000000000000000000000000000
00000000000000000000000000000000

0
 000000000000000100100010010100
                               1

*/